LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_arith.all;
USE IEEE.std_logic_signed.all;
use work.adder_Package.all;

PACKAGE OUTPUT_NODE_PACKAGE IS

COMPONENT OUTPUT_NODE
      PORT (x: IN INPUTARRAY;
            clk, rst: IN STD_LOGIC;
            y: OUT INTEGER);
end component;

end package;

-----------------------------------
----------NODE---------------------
-----------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
USE IEEE.std_logic_signed.all;
use work.NODE_Package.all;
use work.MAC_Package.all;
use work.adder_package.all;
use work.LUT_package.all;
use work.OUTPUT_NODE_PACKAGE.all;

entity OUTPUT_NODE is
      PORT (x: IN INPUTARRAY;
      clk, rst: IN STD_LOGIC;
      y: OUT INTEGER);
end OUTPUT_NODE;

architecture NN of OUTPUT_NODE is

SIGNAL output_number : SIGNED(3 DOWNTO 0);
SIGNAL output_value : INTEGER;

begin
    
y <= output_value;

    PROCESS (x,clk)
    BEGIN
        output_number <= x(0);
        for i in 0 to K-1 loop
            IF(x(i) > output_number) THEN
                output_number <= x(i);
                output_value <= i;
            END IF;
        end loop;
    END PROCESS;

end NN;