library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY multiplier  IS 
	PORT( a,  b:  IN  STD_LOGIC_VECTOR  (3  DOWNTO  0);       
		  prod:  OUT  STD_LOGIC_VECTOR  (7  DOWNTO  0)); 
END multiplier; 

architecture dataflow of multiplier is

begin

end architecture ; -- dataflow